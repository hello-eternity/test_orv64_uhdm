`define PYGMY_ES1Y
