
module or_gate # (
  parameter WIDTH = 1
) (
  input   logic [WIDTH-1:0] in_0,
  input   logic [WIDTH-1:0] in_1,
  output  logic [WIDTH-1:0] out
  );

  assign out = in_0 | in_1;

endmodule

module or_gate_24 # (
  parameter WIDTH = 1
) (
  input   logic [WIDTH-1:0] in_0,
  input   logic [WIDTH-1:0] in_1,
  input   logic [WIDTH-1:0] in_2,
  input   logic [WIDTH-1:0] in_3,
  input   logic [WIDTH-1:0] in_4,
  input   logic [WIDTH-1:0] in_5,
  input   logic [WIDTH-1:0] in_6,
  input   logic [WIDTH-1:0] in_7,
  input   logic [WIDTH-1:0] in_8,
  input   logic [WIDTH-1:0] in_9,
  input   logic [WIDTH-1:0] in_10,
  input   logic [WIDTH-1:0] in_11,
  input   logic [WIDTH-1:0] in_12,
  input   logic [WIDTH-1:0] in_13,
  input   logic [WIDTH-1:0] in_14,
  input   logic [WIDTH-1:0] in_15,
  input   logic [WIDTH-1:0] in_16,
  input   logic [WIDTH-1:0] in_17,
  input   logic [WIDTH-1:0] in_18,
  input   logic [WIDTH-1:0] in_19,
  input   logic [WIDTH-1:0] in_20,
  input   logic [WIDTH-1:0] in_21,
  input   logic [WIDTH-1:0] in_22,
  input   logic [WIDTH-1:0] in_23,
  output  logic [WIDTH-1:0] out
  );

  assign out = in_0 | in_1 | in_2 | in_3 | in_4 | in_5 | in_6 | in_7 | in_8 | in_9 | in_10 | in_11 | in_12 | in_13 | in_14 | in_15 | in_16 | in_17 | in_18 | in_19 | in_20 | in_21 | in_22 | in_23;

endmodule

