`define FPGA
`define SYNTHESIS
`define ORV64_SUPPORT_MULDIV
`define ORV64_SUPPORT_HPMCOUNTER
